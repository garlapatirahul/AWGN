module square_root_coeff (
    
    input clk,                    // system clock
 
    // Data interface
    input [5:0] addr,             // read address
    output reg [19:0] c0,         // coefficient c0, 
    output reg [11:0] c1,         // coefficient c1, 
              
);
 
// Local variables
reg [30:0] d;    // {c0, c1}
 
 
// Table
always @ (*) begin
    case (addr)
        8'd0  : d = 32'b1100110111110001110_011110000000;
        8'd1  : d = 32'b1101001011111011001_111011110011;
        8'd2  : d = 32'b0101010111101101110_010101000000;
        8'd3  : d = 32'b1101011101111111001_111111010011;
        8'd4  : d = 32'b0101100101100100010_101110011100;
        8'd5  : d = 32'b1101111010111110111_101000001100;
        8'd6  : d = 32'b1110001001011101011_011011010011;
        8'd7  : d = 32'b1110010011110011100_101101011001;
        8'd8  : d = 32'b0101111110110101010_011001000110;
        8'd9  : d = 32'b1110010010111100001_111010111011;
        8'd10 : d = 32'b0110100000101110001_000111111000;
        8'd11 : d = 32'b0110101010110001001_101100100011;
        8'd12 : d = 32'b0110001111001100101_111001100011;
        8'd13 : d = 32'b1110100001110101001_111010010101;
        8'd14 : d = 32'b0110101110100111010_011010000101;
        8'd15 : d = 32'b1110110111111100110_001011001010;
        8'd16 : d = 32'b0110011010110100101_100100110110;
        8'd17 : d = 32'b0110101100001001100_111111010010;
        8'd18 : d = 32'b0110111000000001000_101110011111;
        8'd19 : d = 32'b11111000000101011011_101001101001;
        8'd20 : d = 32'b00110100011100101111_011100100011;
        8'd21 : d = 32'b00110110011110011100_001100101001;
        8'd22 : d = 32'b10110111110111000110_001000110100;
        8'd23 : d = 32'b00111000110111101101_001100011100;
        8'd24 : d = 32'b10110101010011111110_011110111110;
        8'd25 : d = 32'b00110111001110000100_100001100011;
        8'd26 : d = 32'b00111000100001011001_101000110010;
        8'd27 : d = 32'b11111001011110000001_110011100100;
        8'd28 : d = 32'b01110110000000110101_101010001000;
        8'd29 : d = 32'b11110111110100011001_111100101010;
        8'd30 : d = 32'b11111001000011001010_001101011010;
        8'd31 : d = 32'b10111001111100011001_011110010110;
        8'd32 : d = 32'b01110110100110001001_111100010101;
        8'd33 : d = 32'b11111000010100000101_011100110010;
        8'd34 : d = 32'b10111001011110111001_110101110100;
        8'd35 : d = 32'b11111010010101001100_001100000110;
        8'd36 : d = 32'b00110111000101110100_010100010001;
        8'd37 : d = 32'b01111000101110110010_000000111110;
        8'd38 : d = 32'b10111001110110001010_100001010001;
        8'd39 : d = 32'b10111010101001111011_111100001111;
        8'd40 : d = 32'b00110111100001000101_110000110111;
        8'd41 : d = 32'b11111001000101101101_101000011110;
        8'd42 : d = 32'b11111010001010000011_001111001101;
        8'd43 : d = 32'b00111010111011100011_101110010101;
        8'd44 : d = 32'b01110111111000111001_010001010110;
        8'd45 : d = 32'b00111001011001101000_010010101101;
        8'd46 : d = 32'b01111010011011010001_111111001101;
        8'd47 : d = 32'b11111011001010110011_100010000001;
        8'd48 : d = 32'b01111000001101111010_110101000100;
        8'd49 : d = 32'b11111001101011001001_111111001110;
        8'd50 : d = 32'b00111010101010011000_110000111001;
        8'd51 : d = 32'b11111011011000001000_010111000010;
        8'd52 : d = 32'b11111000100000100111_011011100010;
        8'd53 : d = 32'b11111001111010101101_101101101001;
        8'd54 : d = 32'b01111010110111110001_100100000001;
        8'd55 : d = 32'b01111011100011111010_001101001010;
        8'd56 : d = 32'b10111000110001011010_000100010101;
        8'd57 : d = 32'b00111010001000101001_011101101101;
        8'd58 : d = 32'b00111011000011101110_011000010110;
        8'd59 : d = 32'b10111011101110011011_000100001110;
        8'd60 : d = 32'b11111001000000100110_101111001000;
        8'd61 : d = 32'b01111010010101001110_001111001011;
        8'd62 : d = 32'b01111011001110100000_001101101110;
        8'd63 : d = 32'b11111011110111111001_111100000110;
        default: d = 31'd0;
    endcase
end
 
 
// Output data
always @ (posedge clk) begin
    c0 <= d[31:12];
    c1 <= d[11:0];
end
 
 
endmodule
