
module sin_cos_coeff (
    
    input clk,                    // system clock
 
    // Data interface
    input [6:0] addr,             // read address
    output reg [18:0] c0,         // coefficient c0, 
    output reg [11:0] c1,         // coefficient c1, 
              
);
 
// Local variables
reg [30:0] d;    // {c0, c1}
 
 
// Table
always @ (*) begin
    case (addr)
        8'd0  : d = 31'b1100110111110001110_011110000000;
        8'd1  : d = 31'b1101001011111011001_111011110011;
        8'd2  : d = 31'b0101010111101101110_010101000000;
        8'd3  : d = 31'b1101011101111111001_111111010011;
        8'd4  : d = 31'b0101100101100100010_101110011100;
        8'd5  : d = 31'b1101111010111110111_101000001100;
        8'd6  : d = 31'b1110001001011101011_011011010011;
        8'd7  : d = 31'b1110010011110011100_101101011001;
        8'd8  : d = 31'b0101111110110101010_011001000110;
        8'd9  : d = 31'b1110010010111100001_111010111011;
        8'd10 : d = 31'b0110100000101110001_000111111000;
        8'd11 : d = 31'b0110101010110001001_101100100011;
        8'd12 : d = 31'b0110001111001100101_111001100011;
        8'd13 : d = 31'b1110100001110101001_111010010101;
        8'd14 : d = 31'b0110101110100111010_011010000101;
        8'd15 : d = 31'b1110110111111100110_001011001010;
        8'd16 : d = 31'b0110011010110100101_100100110110;
        8'd17 : d = 31'b0110101100001001100_111111010010;
        8'd18 : d = 31'b0110111000000001000_101110011111;
        8'd19 : d = 31'b000111101011110111_111000000101011011_101001101001;
        8'd20 : d = 31'b001001101010111000_110100011100101111_011100100011;
        8'd21 : d = 31'b001001010101110100_110110011110011100_001100101001;
        8'd22 : d = 31'b001001000100001010_110111110111000110_001000110100;
        8'd23 : d = 31'b001000110100111000_111000110111101101_001100011100;
        8'd24 : d = 31'b001010101000111110_110101010011111110_011110111110;
        8'd25 : d = 31'b001010010101100000_110111001110000100_100001100011;
        8'd26 : d = 31'b001010000101010000_111000100001011001_101000110010;
        8'd27 : d = 31'b001001110111001111_111001011110000001_110011100100;
        8'd28 : d = 31'b001011100010101101_110110000000110101_101010001000;
        8'd29 : d = 31'b001011010000100011_110111110100011001_111100101010;
        8'd30 : d = 31'b001011000001011011_111001000011001010_001101011010;
        8'd31 : d = 31'b001010110100011010_111001111100011001_011110010110;
        8'd32 : d = 31'b001100011000111001_110110100110001001_111100010101;
        8'd33 : d = 31'b001100000111110011_111000010100000101_011100110010;
        8'd34 : d = 31'b001011111001100110_111001011110111001_110101110100;
        8'd35 : d = 31'b001011101101011011_111010010101001100_001100000110;
        8'd36 : d = 31'b001101001100000100_110111000101110100_010100010001;
        8'd37 : d = 31'b001100111011111001_111000101110110010_000000111110;
        8'd38 : d = 31'b001100101110011110_111001110110001010_100001010001;
        8'd39 : d = 31'b001100100010111110_111010101001111011_111100001111;
        8'd40 : d = 31'b001101111100101100_110111100001000101_110000110111;
        8'd41 : d = 31'b001101101101010011_111001000101101101_101000011110;
        8'd42 : d = 31'b001101100000100011_111010001010000011_001111001101;
        8'd43 : d = 31'b001101010101101000_111010111011100011_101110010101;
        8'd44 : d = 31'b001110101011000101_110111111000111001_010001010110;
        8'd45 : d = 31'b001110011100011000_111001011001101000_010010101101;
        8'd46 : d = 31'b001110010000001101_111010011011010001_111111001101;
        8'd47 : d = 31'b001110000101110011_111011001010110011_100010000001;
        8'd48 : d = 31'b001111010111100001_111000001101111010_110101000100;
        8'd49 : d = 31'b001111001001011011_111001101011001001_111111001110;
        8'd50 : d = 31'b001110111101110000_111010101010011000_110000111001;
        8'd51 : d = 31'b001110110011110011_111011011000001000_010111000010;
        8'd52 : d = 31'b010000000010001111_111000100000100111_011011100010;
        8'd53 : d = 31'b001111110100101011_111001111010101101_101101101001;
        8'd54 : d = 31'b001111101001011101_111010110111110001_100100000001;
        8'd55 : d = 31'b001111011111111001_111011100011111010_001101001010;
        8'd56 : d = 31'b010000101011011010_111000110001011010_000100010101;
        8'd57 : d = 31'b010000011110010100_111010001000101001_011101101101;
        8'd58 : d = 31'b010000010011100000_111011000011101110_011000010110;
        8'd59 : d = 31'b010000001010010010_111011101110011011_000100001110;
        8'd60 : d = 31'b010001010011001011_111001000000100110_101111001000;
        8'd61 : d = 31'b010001000110100001_111010010101001110_001111001011;
        8'd62 : d = 31'b010000111100000101_111011001110100000_001101101110;
        8'd63 : d = 31'b010000110011001011_111011110111111001_111100000110;
        8'd64 : d = 31'b010001111001101011_111001001110011010_011011101011;
        8'd65 : d = 31'b010001101101011010_111010100000101000_000001110110;
        8'd66 : d = 31'b010001100011010011_111011011000010001_000011111111;
        8'd67 : d = 31'b010001011010101100_111100000000011100_110100101010;
        8'd68 : d = 31'b010010011111000010_111001011011000010_001001101111;
        8'd69 : d = 31'b010010010011001000_111010101011000011_110101100101;
        8'd70 : d = 31'b010010001001010100_111011100001001011_111011000011;
        8'd71 : d = 31'b010010000000111110_111100001000001111_101101110101;
        8'd72 : d = 31'b010011000011010100_111001100110101010_111001001001;
        8'd73 : d = 31'b010010110111110000_111010110100101000_101010001111;
        8'd74 : d = 31'b010010101110001110_111011101001010101_110010110010;
        8'd75 : d = 31'b010010100110000111_111100001111011000_100111100001;
        8'd76 : d = 31'b010011100110101001_111001110001011000_101001101110;
        8'd77 : d = 31'b010011011011011000_111010111101011100_011111101110;
        8'd78 : d = 31'b010011010010000110_111011110000110110_101011000111;
        8'd79 : d = 31'b010011001010001101_111100010101111100_100001101100;
        8'd80 : d = 31'b010100001001000100_111001111011010100_011011010110;
        8'd81 : d = 31'b010011111110000101_111011000101100111_010101111010;
        8'd82 : d = 31'b010011110101000010_111011110111110011_100011111111;
        8'd83 : d = 31'b010011101101010110_111100011100000001_011100010000;
        8'd84 : d = 31'b010100101010101001_111010000100100011_001101111010;
        8'd85 : d = 31'b010100011111111011_111011001101001100_001100110000;
        8'd86 : d = 31'b010100010111000110_111011111110010000_011101010101;
        8'd87 : d = 31'b010100001111100110_111100100001101001_010111001100;
        8'd88 : d = 31'b010101001011011100_111010001101001011_000001010100;
        8'd89 : d = 31'b010101000000111110_111011010100010000_000100001100;
        8'd90 : d = 31'b010100111000010110_111100000100010001_010111000110;
        8'd91 : d = 31'b010100110001000001_111100100110111000_10010011100;
        8'd92 : d = 31'b010101101011100000_111010010101001111_110101011110;
        8'd93 : d = 31'b010101100001010001_111011011010111000_111100001000;
        8'd94 : d = 31'b010101011000110110_111100001001111000_010001010000;
        8'd95 : d = 31'b010101010001101011_111100101011110001_001110000000;
        8'd96 : d = 31'b010110001010111001_111010011100110100_101010010101;
        8'd97 : d = 31'b010110000000110111_111011100001000100_110100100011;
        8'd98 : d = 31'b010101111000101000_111100001111001001_001011110000;
        8'd99 : d = 31'b010101110001100111_111100110000010110_001001110100;
        8'd100: d = 31'b010110101001101001_111010100011111100_011111110011;
        8'd101: d = 31'b010110011111110100_111011100110111001_101101011001;
        8'd102: d = 31'b010110010111101111_111100010100000101_000110100100;
        8'd103: d = 31'b010110010000111000_111100110100101001_000101111000;
        8'd104: d = 31'b010111000111110010_111010101010101010_010101110101;
        8'd105: d = 31'b010110111110001010_111011101100011001_100110101000;
        8'd106: d = 31'b010110110110001111_111100011000101111_000001101010;
        8'd107: d = 31'b010110101111100000_111100111000101100_000010001010;
        8'd108: d = 31'b010111100101010111_111010110001000000_001100011001;
        8'd109: d = 31'b010111011011111010_111011110001100101_100000001110;
        8'd110: d = 31'b010111010100001000_111100011101001000_111101000001;
        8'd111: d = 31'b010111001101100010_111100111100100000_111110101000;
        8'd112: d = 31'b011000000010011001_111010110111000001_000011011011;
        8'd113: d = 31'b010111111001000111_111011110110011111_011010001001;
        8'd114: d = 31'b010111110001011110_111100100001010011_111000100111;
        8'd115: d = 31'b010111101011000000_111101000000000111_111011010010;
        8'd116: d = 31'b011000011110111010_111010111100101110_111010111001;
        8'd117: d = 31'b011000010101110010_111011111011001001_010100010111;
        8'd118: d = 31'b011000001110010011_111100100101001111_110100011011;
        8'd119: d = 31'b011000000111111011_111101000011100010_111000000111;
        8'd120: d = 31'b011000111010111100_111011000010001010_110010110001;
        8'd121: d = 31'b011000110001111110_111011111111100100_001110110111;
        8'd122: d = 31'b011000101010100111_111100101000111110_110000011100;
        8'd123: d = 31'b011000100100010110_111101000110110010_110101000110;
        8'd124: d = 31'b011001010110100001_111011000111010100_101011000001;
        8'd125: d = 31'b011001001101101100_111100000011110001_001001100110;
        8'd126: d = 31'b011001000110011100_111100101100100010_101100101001;
        8'd127: d = 31'b011001000000010011_111101001001111000_110010001110;
        default: d = 31'd0;
    endcase
end
 
 
// Output data
always @ (posedge clk) begin
    c0 <= d[30:12];
    c1 <= d[11:0];
end
 
 
endmodule
