module AWGN(Clock, reset, urng_seed1, urng_seed2, urng_seed3, urng_seed4, urng_seed5, urng_seed6, awgn_out)

input Clock,reset, urng_seed1, urng_seed2, urng_seed3, urng_seed4, urng_seed5, urng_seed6;
output awgn_out;


