
module sin_cos_coeff (
    
    input clk,                    // system clock
 
    // Data interface
    input [6:0] addr,             // read address
    output reg [18:0] c0,         // coefficient c0, 
    output reg [11:0] c1,         // coefficient c1, 
              
);
 
// Local variables
reg [30:0] d;    // {c0, c1}
 
 
// Table
always @ (*) begin
    case (addr)
        8'd0  : d = 31'b1100110111110001110_011110000000;
        8'd1  : d = 31'b1101001011111011001_111011110011;
        8'd2  : d = 31'b0101010111101101110_010101000000;
        8'd3  : d = 31'b1101011101111111001_111111010011;
        8'd4  : d = 31'b0101100101100100010_101110011100;
        8'd5  : d = 31'b1101111010111110111_101000001100;
        8'd6  : d = 31'b1110001001011101011_011011010011;
        8'd7  : d = 31'b1110010011110011100_101101011001;
        8'd8  : d = 31'b0101111110110101010_011001000110;
        8'd9  : d = 31'b1110010010111100001_111010111011;
        8'd10 : d = 31'b0110100000101110001_000111111000;
        8'd11 : d = 31'b0110101010110001001_101100100011;
        8'd12 : d = 31'b0110001111001100101_111001100011;
        8'd13 : d = 31'b1110100001110101001_111010010101;
        8'd14 : d = 31'b0110101110100111010_011010000101;
        8'd15 : d = 31'b1110110111111100110_001011001010;
        8'd16 : d = 31'b0110011010110100101_100100110110;
        8'd17 : d = 31'b0110101100001001100_111111010010;
        8'd18 : d = 31'b0110111000000001000_101110011111;
        8'd19 : d = 31'b0001111010111101111_101001101001;
        8'd20 : d = 31'b0010011010101110001_011100100011;
        8'd21 : d = 31'b0010010101011101001_001100101001;
        8'd22 : d = 31'b0010010001000010101_001000110100;
        8'd23 : d = 31'b0010001101001110001_001100011100;
        8'd24 : d = 31'b0010101010001111101_011110111110;
        8'd25 : d = 31'b0010100101011000001_100001100011;
        8'd26 : d = 31'b0010100001010100001_101000110010;
        8'd27 : d = 31'b0010011101110011111_110011100100;
        8'd28 : d = 31'b0010111000101011011_101010001000;
        8'd29 : d = 31'b0010110100001000111_111100101010;
        8'd30 : d = 31'b0010110000010110111_001101011010;
        8'd31 : d = 31'b0010101101000110101_011110010110;
        8'd32 : d = 31'b0011000110001110011_111100010101;
        8'd33 : d = 31'b0011000001111100111_011100110010;
        8'd34 : d = 31'b0010111110011001101_110101110100;
        8'd35 : d = 31'b0010111011010110111_001100000110;
        8'd36 : d = 31'b0011010011000001001_010100010001;
        8'd37 : d = 31'b0011001110111110011_000000111110;
        8'd38 : d = 31'b0011001011100111101_100001010001;
        8'd39 : d = 31'b0011001000101111101_111100001111;
        8'd40 : d = 31'b0011011111001011001_110000110111;
        8'd41 : d = 31'b0011011011010100111_101000011110;
        8'd42 : d = 31'b0011011000001000111_001111001101;
        8'd43 : d = 31'b0011010101011010001_101110010101;
        8'd44 : d = 31'b0011101010110001011_010001010110;
        8'd45 : d = 31'b0011100111000110001_010010101101;
        8'd46 : d = 31'b0011100100000011011_111111001101;
        8'd47 : d = 31'b0011100001011100111_100010000001;
        8'd48 : d = 31'b0011110101111000011_110101000100;
        8'd49 : d = 31'b0011110010010110111_111111001110;
        8'd50 : d = 31'b0011101111011100001_110000111001;
        8'd51 : d = 31'b0011101100111100111_010111000010;
        8'd52 : d = 31'b0100000000100011111_011011100010;
        8'd53 : d = 31'b0011111101001010111_101101101001;
        8'd54 : d = 31'b0011111010010111011_100100000001;
        8'd55 : d = 31'b0011110111111110011_001101001010;
        8'd56 : d = 31'b0100001010110110101_000100010101;
        8'd57 : d = 31'b0100000111100101001_011101101101;
        8'd58 : d = 31'b0100000100111000001_011000010110;
        8'd59 : d = 31'b0100000010100100101_000100001110;
        8'd60 : d = 31'b0100010100110010111_101111001000;
        8'd61 : d = 31'b0100010001101000011_001111001011;
        8'd62 : d = 31'b0100001111000001011_001101101110;
        8'd63 : d = 31'b0100001100110010111_111100000110;
        8'd64 : d = 31'b0100011110011010111_011011101011;
        8'd65 : d = 31'b0100011011010110101_000001110110;
        8'd66 : d = 31'b0100011000110100111_000011111111;
        8'd67 : d = 31'b0100010110101011001_110100101010;
        8'd68 : d = 31'b0100100111110000101_001001101111;
        8'd69 : d = 31'b0100100100110010001_110101100101;
        8'd70 : d = 31'b0100100010010101001_111011000011;
        8'd71 : d = 31'b0100100000001111101_101101110101;
        8'd72 : d = 31'b0100110000110101001_111001001001;
        8'd73 : d = 31'b0100101101111100001_101010001111;
        8'd74 : d = 31'b0100101011100011101_110010110010;
        8'd75 : d = 31'b0100101001100001111_100111100001;
        8'd76 : d = 31'b0100111001101010011_101001101110;
        8'd77 : d = 31'b0100110110110110001_011111101110;
        8'd78 : d = 31'b0100110100100001101_101011000111;
        8'd79 : d = 31'b0100110010100011011_100001101100;
        8'd80 : d = 31'b0101000010010001001_011011010110;
        8'd81 : d = 31'b0100111111100001011_010101111010;
        8'd82 : d = 31'b0100111101010000101_100011111111;
        8'd83 : d = 31'b0100111011010101101_011100010000;
        8'd84 : d = 31'b0101001010101010011_001101111010;
        8'd85 : d = 31'b0101000111111110111_001100110000;
        8'd86 : d = 31'b0101000101110001101_011101010101;
        8'd87 : d = 31'b0101000011111001101_010111001100;
        8'd88 : d = 31'b0101010010110111001_000001010100;
        8'd89 : d = 31'b0101010000001111101_000100001100;
        8'd90 : d = 31'b0101001110000101101_010111000110;
        8'd91 : d = 31'b0101001100010000011_10010011100;
        8'd92 : d = 31'b0101011010111000001_110101011110;
        8'd93 : d = 31'b0101011000010100011_111100001000;
        8'd94 : d = 31'b0101010110001101101_010001010000;
        8'd95 : d = 31'b0101010100011010111_001110000000;
        8'd96 : d = 31'b0101100010101110011_101010010101;
        8'd97 : d = 31'b0101100000001101111_110100100011;
        8'd98 : d = 31'b0101011110001010001_001011110000;
        8'd99 : d = 31'b0101011100011001111_001001110100;
        8'd100: d = 31'b0101101010011010011_011111110011;
        8'd101: d = 31'b0101100111111101001_101101011001;
        8'd102: d = 31'b0101100101111011111_000110100100;
        8'd103: d = 31'b0101100100001110001_000101111000;
        8'd104: d = 31'b0101110001111100101_010101110101;
        8'd105: d = 31'b0101101111100010101_100110101000;
        8'd106: d = 31'b0101101101100011111_000001101010;
        8'd107: d = 31'b0101101011111000001_000010001010;
        8'd108: d = 31'b0101111001010101111_001100011001;
        8'd109: d = 31'b0101110110111110101_100000001110;
        8'd110: d = 31'b0101110101000010001_111101000001;
        8'd111: d = 31'b0101110011011000101_111110101000;
        8'd112: d = 31'b0110000000100110011_000011011011;
        8'd113: d = 31'b0101111110010001111_011010001001;
        8'd114: d = 31'b0101111100010111101_111000100111;
        8'd115: d = 31'b0101111010110000001_111011010010;
        8'd116: d = 31'b0110000111101110101_111010111001;
        8'd117: d = 31'b0110000101011100101_010100010111;
        8'd118: d = 31'b0110000011100100111_110100011011;
        8'd119: d = 31'b0110000001111110111_111000000111;
        8'd120: d = 31'b0110001110101111001_110010110001;
        8'd121: d = 31'b0110001100011111101_001110110111;
        8'd122: d = 31'b0110001010101001111_110000011100;
        8'd123: d = 31'b0110001001000101101_110101000110;
        8'd124: d = 31'b0110010101101000011_101011000001;
        8'd125: d = 31'b0110010011011011001_001001100110;
        8'd126: d = 31'b0110010001100111001_101100101001;
        8'd127: d = 31'b0110010000000100111_110010001110;
        default: d = 31'd0;
    endcase
end
 
 
// Output data
always @ (posedge clk) begin
    c0 <= d[30:12];
    c1 <= d[11:0];
end
 
 
endmodule
